-- megafunction wizard: %Parallel Flash Loader%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altparallel_flash_loader 

-- ============================================================
-- File Name: p2.vhd
-- Megafunction Name(s):
-- 			altparallel_flash_loader
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.1 Build 646 04/11/2019 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2019  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY p2 IS
	PORT
	(
		fpga_conf_done		: IN STD_LOGIC ;
		fpga_nstatus		: IN STD_LOGIC ;
		fpga_pgm		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		pfl_clk		: IN STD_LOGIC ;
		pfl_flash_access_granted		: IN STD_LOGIC ;
		pfl_nreconfigure		: IN STD_LOGIC  := '1';
		pfl_nreset		: IN STD_LOGIC ;
		flash_addr		: OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
		flash_clk		: OUT STD_LOGIC ;
		flash_data		: INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		flash_nadv		: OUT STD_LOGIC ;
		flash_nce		: OUT STD_LOGIC ;
		flash_noe		: OUT STD_LOGIC ;
		flash_nreset		: OUT STD_LOGIC ;
		flash_nwe		: OUT STD_LOGIC ;
		fpga_data		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		fpga_dclk		: OUT STD_LOGIC ;
		fpga_nconfig		: OUT STD_LOGIC ;
		pfl_flash_access_request		: OUT STD_LOGIC 
	);
END p2;


ARCHITECTURE SYN OF p2 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (24 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC ;
	SIGNAL sub_wire3	: STD_LOGIC ;
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC ;
	SIGNAL sub_wire6	: STD_LOGIC ;
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC ;
	SIGNAL sub_wire9	: STD_LOGIC ;
	SIGNAL sub_wire10	: STD_LOGIC ;



	COMPONENT altparallel_flash_loader
	GENERIC (
		addr_width		: NATURAL;
		burst_mode		: NATURAL;
		burst_mode_intel		: NATURAL;
		burst_mode_latency_count		: NATURAL;
		burst_mode_numonyx		: NATURAL;
		burst_mode_spansion		: NATURAL;
		clk_divisor		: NATURAL;
		conf_data_width		: NATURAL;
		conf_wait_timer_width		: NATURAL;
		dclk_divisor		: NATURAL;
		decompressor_mode		: STRING;
		features_cfg		: NATURAL;
		features_pgm		: NATURAL;
		flash_burst_extra_cycle		: NATURAL;
		flash_data_width		: NATURAL;
		flash_nreset_checkbox		: NATURAL;
		flash_nreset_counter		: NATURAL;
		flash_type		: STRING;
		normal_mode		: NATURAL;
		n_flash		: NATURAL;
		option_bits_start_address		: NATURAL;
		page_clk_divisor		: NATURAL;
		page_mode		: NATURAL;
		qspi_data_delay		: NATURAL;
		qspi_data_delay_count		: NATURAL;
		safe_mode_halt		: NATURAL;
		safe_mode_retry		: NATURAL;
		safe_mode_revert		: NATURAL;
		safe_mode_revert_addr		: NATURAL;
		tristate_checkbox		: NATURAL;
		lpm_type		: STRING
	);
	PORT (
			fpga_conf_done	: IN STD_LOGIC ;
			fpga_nstatus	: IN STD_LOGIC ;
			fpga_pgm	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			pfl_clk	: IN STD_LOGIC ;
			pfl_flash_access_granted	: IN STD_LOGIC ;
			pfl_nreconfigure	: IN STD_LOGIC ;
			pfl_nreset	: IN STD_LOGIC ;
			flash_addr	: OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
			flash_clk	: OUT STD_LOGIC ;
			flash_nadv	: OUT STD_LOGIC ;
			flash_nce	: OUT STD_LOGIC ;
			flash_noe	: OUT STD_LOGIC ;
			flash_nreset	: OUT STD_LOGIC ;
			flash_nwe	: OUT STD_LOGIC ;
			fpga_data	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			fpga_dclk	: OUT STD_LOGIC ;
			fpga_nconfig	: OUT STD_LOGIC ;
			pfl_flash_access_request	: OUT STD_LOGIC ;
			flash_data	: INOUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	flash_addr    <= sub_wire0(24 DOWNTO 0);
	flash_clk    <= sub_wire1;
	flash_nadv    <= sub_wire2;
	flash_nce    <= sub_wire3;
	flash_noe    <= sub_wire4;
	flash_nreset    <= sub_wire5;
	flash_nwe    <= sub_wire6;
	fpga_data    <= sub_wire7(15 DOWNTO 0);
	fpga_dclk    <= sub_wire8;
	fpga_nconfig    <= sub_wire9;
	pfl_flash_access_request    <= sub_wire10;

	altparallel_flash_loader_component : altparallel_flash_loader
	GENERIC MAP (
		addr_width => 25,
		burst_mode => 1,
		burst_mode_intel => 1,
		burst_mode_latency_count => 3,
		burst_mode_numonyx => 0,
		burst_mode_spansion => 0,
		clk_divisor => 4,
		conf_data_width => 16,
		conf_wait_timer_width => 19,
		dclk_divisor => 1,
		decompressor_mode => "NONE",
		features_cfg => 1,
		features_pgm => 0,
		flash_burst_extra_cycle => 0,
		flash_data_width => 16,
		flash_nreset_checkbox => 0,
		flash_nreset_counter => 2500,
		flash_type => "CFI_FLASH",
		normal_mode => 0,
		n_flash => 1,
		option_bits_start_address => 98304,
		page_clk_divisor => 1,
		page_mode => 0,
		qspi_data_delay => 0,
		qspi_data_delay_count => 1,
		safe_mode_halt => 0,
		safe_mode_retry => 1,
		safe_mode_revert => 0,
		safe_mode_revert_addr => 0,
		tristate_checkbox => 1,
		lpm_type => "altparallel_flash_loader"
	)
	PORT MAP (
		fpga_conf_done => fpga_conf_done,
		fpga_nstatus => fpga_nstatus,
		fpga_pgm => fpga_pgm,
		pfl_clk => pfl_clk,
		pfl_flash_access_granted => pfl_flash_access_granted,
		pfl_nreconfigure => pfl_nreconfigure,
		pfl_nreset => pfl_nreset,
		flash_addr => sub_wire0,
		flash_clk => sub_wire1,
		flash_nadv => sub_wire2,
		flash_nce => sub_wire3,
		flash_noe => sub_wire4,
		flash_nreset => sub_wire5,
		flash_nwe => sub_wire6,
		fpga_data => sub_wire7,
		fpga_dclk => sub_wire8,
		fpga_nconfig => sub_wire9,
		pfl_flash_access_request => sub_wire10,
		flash_data => flash_data
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: CLOCK_FREQUENCY_EDIT STRING "50"
-- Retrieval info: PRIVATE: DCLK_DIVISOR_COMBO STRING "1"
-- Retrieval info: PRIVATE: FLASH_ACCESS_TIME_EDIT STRING "100"
-- Retrieval info: PRIVATE: IDC_DECOMPRESSOR_COMBO STRING "None"
-- Retrieval info: PRIVATE: IDC_FLASH_DATA_WIDTH_COMBO STRING "16 bits"
-- Retrieval info: PRIVATE: IDC_FLASH_DEVICE_COMBO STRING "CFI 512 Mbit"
-- Retrieval info: PRIVATE: IDC_FLASH_NRESET_CHECKBOX STRING "1"
-- Retrieval info: PRIVATE: IDC_FLASH_TYPE_COMBO STRING "CFI Parallel Flash"
-- Retrieval info: PRIVATE: IDC_FPGA_CONF_SCHEME_COMBO STRING "FPP x16 (fast passive parallel x16)"
-- Retrieval info: PRIVATE: IDC_NUM_FLASH_COMBO STRING "1"
-- Retrieval info: PRIVATE: IDC_OPERATING_MODES_COMBO STRING "FPGA Configuration"
-- Retrieval info: PRIVATE: IDC_READ_MODES_COMBO STRING "Intel Burst Mode with 3 LC (P30 or P33 only)"
-- Retrieval info: PRIVATE: IDC_SAFE_MODE_COMBO STRING "Retry same page"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX V"
-- Retrieval info: PRIVATE: OPTION_BIT_ADDRESS_EDIT STRING "18000"
-- Retrieval info: PRIVATE: RECONFIGURE_CHECKBOX STRING "1"
-- Retrieval info: PRIVATE: RSU_WATCHHDOG_CHECKBOX STRING "0"
-- Retrieval info: PRIVATE: RSU_WATCHHDOG_COUNTER_EDIT STRING "100"
-- Retrieval info: PRIVATE: SAFE_MODE_REVERT_EDIT STRING ""
-- Retrieval info: PRIVATE: TRISTATE_CHECKBOX STRING "1"
-- Retrieval info: CONSTANT: ADDR_WIDTH NUMERIC "25"
-- Retrieval info: CONSTANT: BURST_MODE NUMERIC "1"
-- Retrieval info: CONSTANT: BURST_MODE_INTEL NUMERIC "1"
-- Retrieval info: CONSTANT: BURST_MODE_LATENCY_COUNT NUMERIC "3"
-- Retrieval info: CONSTANT: BURST_MODE_NUMONYX NUMERIC "0"
-- Retrieval info: CONSTANT: BURST_MODE_SPANSION NUMERIC "0"
-- Retrieval info: CONSTANT: CLK_DIVISOR NUMERIC "4"
-- Retrieval info: CONSTANT: CONF_DATA_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: CONF_WAIT_TIMER_WIDTH NUMERIC "19"
-- Retrieval info: CONSTANT: DCLK_DIVISOR NUMERIC "1"
-- Retrieval info: CONSTANT: DECOMPRESSOR_MODE STRING "NONE"
-- Retrieval info: CONSTANT: FEATURES_CFG NUMERIC "1"
-- Retrieval info: CONSTANT: FEATURES_PGM NUMERIC "0"
-- Retrieval info: CONSTANT: FLASH_BURST_EXTRA_CYCLE NUMERIC "0"
-- Retrieval info: CONSTANT: FLASH_DATA_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: FLASH_NRESET_CHECKBOX NUMERIC "0"
-- Retrieval info: CONSTANT: FLASH_NRESET_COUNTER NUMERIC "2500"
-- Retrieval info: CONSTANT: FLASH_TYPE STRING "CFI_FLASH"
-- Retrieval info: CONSTANT: NORMAL_MODE NUMERIC "0"
-- Retrieval info: CONSTANT: N_FLASH NUMERIC "1"
-- Retrieval info: CONSTANT: OPTION_BITS_START_ADDRESS NUMERIC "98304"
-- Retrieval info: CONSTANT: PAGE_CLK_DIVISOR NUMERIC "1"
-- Retrieval info: CONSTANT: PAGE_MODE NUMERIC "0"
-- Retrieval info: CONSTANT: QSPI_DATA_DELAY NUMERIC "0"
-- Retrieval info: CONSTANT: QSPI_DATA_DELAY_COUNT NUMERIC "1"
-- Retrieval info: CONSTANT: SAFE_MODE_HALT NUMERIC "0"
-- Retrieval info: CONSTANT: SAFE_MODE_RETRY NUMERIC "1"
-- Retrieval info: CONSTANT: SAFE_MODE_REVERT NUMERIC "0"
-- Retrieval info: CONSTANT: SAFE_MODE_REVERT_ADDR NUMERIC "0"
-- Retrieval info: CONSTANT: TRISTATE_CHECKBOX NUMERIC "1"
-- Retrieval info: USED_PORT: flash_addr 0 0 25 0 OUTPUT NODEFVAL "flash_addr[24..0]"
-- Retrieval info: USED_PORT: flash_clk 0 0 0 0 OUTPUT NODEFVAL "flash_clk"
-- Retrieval info: USED_PORT: flash_data 0 0 16 0 BIDIR NODEFVAL "flash_data[15..0]"
-- Retrieval info: USED_PORT: flash_nadv 0 0 0 0 OUTPUT NODEFVAL "flash_nadv"
-- Retrieval info: USED_PORT: flash_nce 0 0 0 0 OUTPUT NODEFVAL "flash_nce"
-- Retrieval info: USED_PORT: flash_noe 0 0 0 0 OUTPUT NODEFVAL "flash_noe"
-- Retrieval info: USED_PORT: flash_nreset 0 0 0 0 OUTPUT NODEFVAL "flash_nreset"
-- Retrieval info: USED_PORT: flash_nwe 0 0 0 0 OUTPUT NODEFVAL "flash_nwe"
-- Retrieval info: USED_PORT: fpga_conf_done 0 0 0 0 INPUT NODEFVAL "fpga_conf_done"
-- Retrieval info: USED_PORT: fpga_data 0 0 16 0 OUTPUT NODEFVAL "fpga_data[15..0]"
-- Retrieval info: USED_PORT: fpga_dclk 0 0 0 0 OUTPUT NODEFVAL "fpga_dclk"
-- Retrieval info: USED_PORT: fpga_nconfig 0 0 0 0 OUTPUT NODEFVAL "fpga_nconfig"
-- Retrieval info: USED_PORT: fpga_nstatus 0 0 0 0 INPUT NODEFVAL "fpga_nstatus"
-- Retrieval info: USED_PORT: fpga_pgm 0 0 3 0 INPUT NODEFVAL "fpga_pgm[2..0]"
-- Retrieval info: USED_PORT: pfl_clk 0 0 0 0 INPUT NODEFVAL "pfl_clk"
-- Retrieval info: USED_PORT: pfl_flash_access_granted 0 0 0 0 INPUT NODEFVAL "pfl_flash_access_granted"
-- Retrieval info: USED_PORT: pfl_flash_access_request 0 0 0 0 OUTPUT NODEFVAL "pfl_flash_access_request"
-- Retrieval info: USED_PORT: pfl_nreconfigure 0 0 0 0 INPUT VCC "pfl_nreconfigure"
-- Retrieval info: USED_PORT: pfl_nreset 0 0 0 0 INPUT NODEFVAL "pfl_nreset"
-- Retrieval info: CONNECT: @fpga_conf_done 0 0 0 0 fpga_conf_done 0 0 0 0
-- Retrieval info: CONNECT: @fpga_nstatus 0 0 0 0 fpga_nstatus 0 0 0 0
-- Retrieval info: CONNECT: @fpga_pgm 0 0 3 0 fpga_pgm 0 0 3 0
-- Retrieval info: CONNECT: @pfl_clk 0 0 0 0 pfl_clk 0 0 0 0
-- Retrieval info: CONNECT: @pfl_flash_access_granted 0 0 0 0 pfl_flash_access_granted 0 0 0 0
-- Retrieval info: CONNECT: @pfl_nreconfigure 0 0 0 0 pfl_nreconfigure 0 0 0 0
-- Retrieval info: CONNECT: @pfl_nreset 0 0 0 0 pfl_nreset 0 0 0 0
-- Retrieval info: CONNECT: flash_addr 0 0 25 0 @flash_addr 0 0 25 0
-- Retrieval info: CONNECT: flash_clk 0 0 0 0 @flash_clk 0 0 0 0
-- Retrieval info: CONNECT: flash_data 0 0 16 0 @flash_data 0 0 16 0
-- Retrieval info: CONNECT: flash_nadv 0 0 0 0 @flash_nadv 0 0 0 0
-- Retrieval info: CONNECT: flash_nce 0 0 0 0 @flash_nce 0 0 0 0
-- Retrieval info: CONNECT: flash_noe 0 0 0 0 @flash_noe 0 0 0 0
-- Retrieval info: CONNECT: flash_nreset 0 0 0 0 @flash_nreset 0 0 0 0
-- Retrieval info: CONNECT: flash_nwe 0 0 0 0 @flash_nwe 0 0 0 0
-- Retrieval info: CONNECT: fpga_data 0 0 16 0 @fpga_data 0 0 16 0
-- Retrieval info: CONNECT: fpga_dclk 0 0 0 0 @fpga_dclk 0 0 0 0
-- Retrieval info: CONNECT: fpga_nconfig 0 0 0 0 @fpga_nconfig 0 0 0 0
-- Retrieval info: CONNECT: pfl_flash_access_request 0 0 0 0 @pfl_flash_access_request 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL p2.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL p2.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL p2.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL p2.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL p2_inst.vhd TRUE
-- Retrieval info: LIB_FILE: altera_mf
