// q_sys.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module q_sys (
		input  wire  clk_clk,                             //                      clk.clk
		inout  wire  opencores_i2c_0_export_0_scl_pad_io, // opencores_i2c_0_export_0.scl_pad_io
		inout  wire  opencores_i2c_0_export_0_sda_pad_io, //                         .sda_pad_io
		input  wire  reset_reset_n,                       //                    reset.reset_n
		input  wire  vj_clk_pls_p_export                  //             vj_clk_pls_p.export
	);

	wire         i2c_cont_bridge_0_avalon_master_chipselect;                   // i2c_cont_bridge_0:mstr_en_n -> mm_interconnect_0:i2c_cont_bridge_0_avalon_master_chipselect
	wire  [31:0] i2c_cont_bridge_0_avalon_master_readdata;                     // mm_interconnect_0:i2c_cont_bridge_0_avalon_master_readdata -> i2c_cont_bridge_0:mstr_data_in
	wire         i2c_cont_bridge_0_avalon_master_waitrequest;                  // mm_interconnect_0:i2c_cont_bridge_0_avalon_master_waitrequest -> i2c_cont_bridge_0:mstr_waitrequest_n
	wire   [9:0] i2c_cont_bridge_0_avalon_master_address;                      // i2c_cont_bridge_0:mstr_address -> mm_interconnect_0:i2c_cont_bridge_0_avalon_master_address
	wire         i2c_cont_bridge_0_avalon_master_read;                         // i2c_cont_bridge_0:mstr_read_n -> mm_interconnect_0:i2c_cont_bridge_0_avalon_master_read
	wire         i2c_cont_bridge_0_avalon_master_write;                        // i2c_cont_bridge_0:mstr_write_n -> mm_interconnect_0:i2c_cont_bridge_0_avalon_master_write
	wire  [31:0] i2c_cont_bridge_0_avalon_master_writedata;                    // i2c_cont_bridge_0:mstr_data_out -> mm_interconnect_0:i2c_cont_bridge_0_avalon_master_writedata
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect;  // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_chipselect -> opencores_i2c_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata;    // opencores_i2c_0:wb_dat_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest; // opencores_i2c_0:wb_ack_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address;     // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_address -> opencores_i2c_0:wb_adr_i
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write;       // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_write -> opencores_i2c_0:wb_we_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata;   // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_writedata -> opencores_i2c_0:wb_dat_i
	wire         vj_avalon_master_0_avalon_master_waitrequest;                 // mm_interconnect_1:vj_avalon_master_0_avalon_master_waitrequest -> vj_avalon_master_0:waitrequest_n
	wire  [31:0] vj_avalon_master_0_avalon_master_readdata;                    // mm_interconnect_1:vj_avalon_master_0_avalon_master_readdata -> vj_avalon_master_0:data_in
	wire         vj_avalon_master_0_avalon_master_read;                        // vj_avalon_master_0:read_n -> mm_interconnect_1:vj_avalon_master_0_avalon_master_read
	wire  [31:0] vj_avalon_master_0_avalon_master_address;                     // vj_avalon_master_0:address -> mm_interconnect_1:vj_avalon_master_0_avalon_master_address
	wire         vj_avalon_master_0_avalon_master_write;                       // vj_avalon_master_0:write_n -> mm_interconnect_1:vj_avalon_master_0_avalon_master_write
	wire  [31:0] vj_avalon_master_0_avalon_master_writedata;                   // vj_avalon_master_0:data_out -> mm_interconnect_1:vj_avalon_master_0_avalon_master_writedata
	wire         mm_interconnect_1_i2c_cont_bridge_0_slv_chipselect;           // mm_interconnect_1:i2c_cont_bridge_0_slv_chipselect -> i2c_cont_bridge_0:slv_en_n
	wire  [31:0] mm_interconnect_1_i2c_cont_bridge_0_slv_readdata;             // i2c_cont_bridge_0:slv_data_out -> mm_interconnect_1:i2c_cont_bridge_0_slv_readdata
	wire         mm_interconnect_1_i2c_cont_bridge_0_slv_waitrequest;          // i2c_cont_bridge_0:slv_waitrequest_n -> mm_interconnect_1:i2c_cont_bridge_0_slv_waitrequest
	wire   [9:0] mm_interconnect_1_i2c_cont_bridge_0_slv_address;              // mm_interconnect_1:i2c_cont_bridge_0_slv_address -> i2c_cont_bridge_0:slv_address
	wire         mm_interconnect_1_i2c_cont_bridge_0_slv_read;                 // mm_interconnect_1:i2c_cont_bridge_0_slv_read -> i2c_cont_bridge_0:slv_read_n
	wire         mm_interconnect_1_i2c_cont_bridge_0_slv_write;                // mm_interconnect_1:i2c_cont_bridge_0_slv_write -> i2c_cont_bridge_0:slv_write_n
	wire  [31:0] mm_interconnect_1_i2c_cont_bridge_0_slv_writedata;            // mm_interconnect_1:i2c_cont_bridge_0_slv_writedata -> i2c_cont_bridge_0:slv_data_in
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [i2c_cont_bridge_0:reset_n, mm_interconnect_0:i2c_cont_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:vj_avalon_master_0_clock_sink_reset_reset_bridge_in_reset_reset, opencores_i2c_0:wb_rst_i, vj_avalon_master_0:reset_n]

	i2c_cont_bridge i2c_cont_bridge_0 (
		.reset_n            (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.clk                (clk_clk),                                             //         clock.clk
		.slv_address        (mm_interconnect_1_i2c_cont_bridge_0_slv_address),     //           slv.address
		.slv_read_n         (~mm_interconnect_1_i2c_cont_bridge_0_slv_read),       //              .read_n
		.slv_write_n        (~mm_interconnect_1_i2c_cont_bridge_0_slv_write),      //              .write_n
		.slv_data_in        (mm_interconnect_1_i2c_cont_bridge_0_slv_writedata),   //              .writedata
		.slv_waitrequest_n  (mm_interconnect_1_i2c_cont_bridge_0_slv_waitrequest), //              .waitrequest_n
		.slv_data_out       (mm_interconnect_1_i2c_cont_bridge_0_slv_readdata),    //              .readdata
		.slv_en_n           (~mm_interconnect_1_i2c_cont_bridge_0_slv_chipselect), //              .chipselect_n
		.mstr_en_n          (i2c_cont_bridge_0_avalon_master_chipselect),          // avalon_master.chipselect_n
		.mstr_address       (i2c_cont_bridge_0_avalon_master_address),             //              .address
		.mstr_write_n       (i2c_cont_bridge_0_avalon_master_write),               //              .write_n
		.mstr_read_n        (i2c_cont_bridge_0_avalon_master_read),                //              .read_n
		.mstr_data_in       (i2c_cont_bridge_0_avalon_master_readdata),            //              .readdata
		.mstr_data_out      (i2c_cont_bridge_0_avalon_master_writedata),           //              .writedata
		.mstr_waitrequest_n (~i2c_cont_bridge_0_avalon_master_waitrequest)         //              .waitrequest_n
	);

	opencores_i2c opencores_i2c_0 (
		.wb_clk_i   (clk_clk),                                                      //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                               //      clock_reset.reset
		.scl_pad_io (opencores_i2c_0_export_0_scl_pad_io),                          //         export_0.export
		.sda_pad_io (opencores_i2c_0_export_0_sda_pad_io),                          //                 .export
		.wb_adr_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  ()                                                              // interrupt_sender.irq
	);

	vj_avalon_master vj_avalon_master_0 (
		.clk           (clk_clk),                                       //       clock_sink.clk
		.reset_n       (~rst_controller_reset_out_reset),               // clock_sink_reset.reset_n
		.read_n        (vj_avalon_master_0_avalon_master_read),         //    avalon_master.read_n
		.write_n       (vj_avalon_master_0_avalon_master_write),        //                 .write_n
		.address       (vj_avalon_master_0_avalon_master_address),      //                 .address
		.data_out      (vj_avalon_master_0_avalon_master_writedata),    //                 .writedata
		.waitrequest_n (~vj_avalon_master_0_avalon_master_waitrequest), //                 .waitrequest_n
		.data_in       (vj_avalon_master_0_avalon_master_readdata),     //                 .readdata
		.clk_pls_p     (vj_clk_pls_p_export)                            //        clk_pls_p.export
	);

	q_sys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                                       //                                     clk_0_clk.clk
		.i2c_cont_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // i2c_cont_bridge_0_reset_reset_bridge_in_reset.reset
		.i2c_cont_bridge_0_avalon_master_address             (i2c_cont_bridge_0_avalon_master_address),                       //               i2c_cont_bridge_0_avalon_master.address
		.i2c_cont_bridge_0_avalon_master_waitrequest         (i2c_cont_bridge_0_avalon_master_waitrequest),                   //                                              .waitrequest
		.i2c_cont_bridge_0_avalon_master_chipselect          (~i2c_cont_bridge_0_avalon_master_chipselect),                   //                                              .chipselect
		.i2c_cont_bridge_0_avalon_master_read                (~i2c_cont_bridge_0_avalon_master_read),                         //                                              .read
		.i2c_cont_bridge_0_avalon_master_readdata            (i2c_cont_bridge_0_avalon_master_readdata),                      //                                              .readdata
		.i2c_cont_bridge_0_avalon_master_write               (~i2c_cont_bridge_0_avalon_master_write),                        //                                              .write
		.i2c_cont_bridge_0_avalon_master_writedata           (i2c_cont_bridge_0_avalon_master_writedata),                     //                                              .writedata
		.opencores_i2c_0_avalon_slave_0_address              (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address),      //                opencores_i2c_0_avalon_slave_0.address
		.opencores_i2c_0_avalon_slave_0_write                (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write),        //                                              .write
		.opencores_i2c_0_avalon_slave_0_readdata             (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata),     //                                              .readdata
		.opencores_i2c_0_avalon_slave_0_writedata            (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata),    //                                              .writedata
		.opencores_i2c_0_avalon_slave_0_waitrequest          (~mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest), //                                              .waitrequest
		.opencores_i2c_0_avalon_slave_0_chipselect           (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect)    //                                              .chipselect
	);

	q_sys_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                                   (clk_clk),                                              //                                                 clk_0_clk.clk
		.vj_avalon_master_0_clock_sink_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // vj_avalon_master_0_clock_sink_reset_reset_bridge_in_reset.reset
		.vj_avalon_master_0_avalon_master_address                        (vj_avalon_master_0_avalon_master_address),             //                          vj_avalon_master_0_avalon_master.address
		.vj_avalon_master_0_avalon_master_waitrequest                    (vj_avalon_master_0_avalon_master_waitrequest),         //                                                          .waitrequest
		.vj_avalon_master_0_avalon_master_read                           (~vj_avalon_master_0_avalon_master_read),               //                                                          .read
		.vj_avalon_master_0_avalon_master_readdata                       (vj_avalon_master_0_avalon_master_readdata),            //                                                          .readdata
		.vj_avalon_master_0_avalon_master_write                          (~vj_avalon_master_0_avalon_master_write),              //                                                          .write
		.vj_avalon_master_0_avalon_master_writedata                      (vj_avalon_master_0_avalon_master_writedata),           //                                                          .writedata
		.i2c_cont_bridge_0_slv_address                                   (mm_interconnect_1_i2c_cont_bridge_0_slv_address),      //                                     i2c_cont_bridge_0_slv.address
		.i2c_cont_bridge_0_slv_write                                     (mm_interconnect_1_i2c_cont_bridge_0_slv_write),        //                                                          .write
		.i2c_cont_bridge_0_slv_read                                      (mm_interconnect_1_i2c_cont_bridge_0_slv_read),         //                                                          .read
		.i2c_cont_bridge_0_slv_readdata                                  (mm_interconnect_1_i2c_cont_bridge_0_slv_readdata),     //                                                          .readdata
		.i2c_cont_bridge_0_slv_writedata                                 (mm_interconnect_1_i2c_cont_bridge_0_slv_writedata),    //                                                          .writedata
		.i2c_cont_bridge_0_slv_waitrequest                               (~mm_interconnect_1_i2c_cont_bridge_0_slv_waitrequest), //                                                          .waitrequest
		.i2c_cont_bridge_0_slv_chipselect                                (mm_interconnect_1_i2c_cont_bridge_0_slv_chipselect)    //                                                          .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
