// q_sys.v

// Generated using ACDS version 12.1sp1 243 at 2013.02.18.13:23:17

`timescale 1 ps / 1 ps
module q_sys (
		inout  wire  opencores_i2c_0_export_0_scl_pad_io, // opencores_i2c_0_export_0.scl_pad_io
		inout  wire  opencores_i2c_0_export_0_sda_pad_io, //                         .sda_pad_io
		input  wire  reset_reset_n,                       //                    reset.reset_n
		input  wire  clk_clk,                             //                      clk.clk
		input  wire  vj_clk_pls_p_export                  //             vj_clk_pls_p.export
	);

	wire         vj_avalon_master_0_avalon_master_waitrequest;                                        // vj_avalon_master_0_avalon_master_translator:av_waitrequest -> vj_avalon_master_0:waitrequest_n
	wire  [31:0] vj_avalon_master_0_avalon_master_writedata;                                          // vj_avalon_master_0:data_out -> vj_avalon_master_0_avalon_master_translator:av_writedata
	wire  [31:0] vj_avalon_master_0_avalon_master_address;                                            // vj_avalon_master_0:address -> vj_avalon_master_0_avalon_master_translator:av_address
	wire         vj_avalon_master_0_avalon_master_write;                                              // vj_avalon_master_0:write_n -> vj_avalon_master_0_avalon_master_translator:av_write
	wire         vj_avalon_master_0_avalon_master_read;                                               // vj_avalon_master_0:read_n -> vj_avalon_master_0_avalon_master_translator:av_read
	wire  [31:0] vj_avalon_master_0_avalon_master_readdata;                                           // vj_avalon_master_0_avalon_master_translator:av_readdata -> vj_avalon_master_0:data_in
	wire         vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_waitrequest;   // i2c_cont_bridge_0_slv_translator:uav_waitrequest -> vj_avalon_master_0_avalon_master_translator:uav_waitrequest
	wire   [2:0] vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_burstcount;    // vj_avalon_master_0_avalon_master_translator:uav_burstcount -> i2c_cont_bridge_0_slv_translator:uav_burstcount
	wire  [31:0] vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_writedata;     // vj_avalon_master_0_avalon_master_translator:uav_writedata -> i2c_cont_bridge_0_slv_translator:uav_writedata
	wire  [31:0] vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_address;       // vj_avalon_master_0_avalon_master_translator:uav_address -> i2c_cont_bridge_0_slv_translator:uav_address
	wire         vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_lock;          // vj_avalon_master_0_avalon_master_translator:uav_lock -> i2c_cont_bridge_0_slv_translator:uav_lock
	wire         vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_write;         // vj_avalon_master_0_avalon_master_translator:uav_write -> i2c_cont_bridge_0_slv_translator:uav_write
	wire         vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_read;          // vj_avalon_master_0_avalon_master_translator:uav_read -> i2c_cont_bridge_0_slv_translator:uav_read
	wire  [31:0] vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdata;      // i2c_cont_bridge_0_slv_translator:uav_readdata -> vj_avalon_master_0_avalon_master_translator:uav_readdata
	wire         vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_debugaccess;   // vj_avalon_master_0_avalon_master_translator:uav_debugaccess -> i2c_cont_bridge_0_slv_translator:uav_debugaccess
	wire   [3:0] vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_byteenable;    // vj_avalon_master_0_avalon_master_translator:uav_byteenable -> i2c_cont_bridge_0_slv_translator:uav_byteenable
	wire         vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdatavalid; // i2c_cont_bridge_0_slv_translator:uav_readdatavalid -> vj_avalon_master_0_avalon_master_translator:uav_readdatavalid
	wire         i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_waitrequest;                    // i2c_cont_bridge_0:slv_waitrequest_n -> i2c_cont_bridge_0_slv_translator:av_waitrequest
	wire  [31:0] i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_writedata;                      // i2c_cont_bridge_0_slv_translator:av_writedata -> i2c_cont_bridge_0:slv_data_in
	wire   [9:0] i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_address;                        // i2c_cont_bridge_0_slv_translator:av_address -> i2c_cont_bridge_0:slv_address
	wire         i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_chipselect;                     // i2c_cont_bridge_0_slv_translator:av_chipselect -> i2c_cont_bridge_0:slv_en_n
	wire         i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_write;                          // i2c_cont_bridge_0_slv_translator:av_write -> i2c_cont_bridge_0:slv_write_n
	wire         i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_read;                           // i2c_cont_bridge_0_slv_translator:av_read -> i2c_cont_bridge_0:slv_read_n
	wire  [31:0] i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_readdata;                       // i2c_cont_bridge_0:slv_data_out -> i2c_cont_bridge_0_slv_translator:av_readdata
	wire         i2c_cont_bridge_0_avalon_master_waitrequest;                                         // i2c_cont_bridge_0_avalon_master_translator:av_waitrequest -> i2c_cont_bridge_0:mstr_waitrequest_n
	wire  [31:0] i2c_cont_bridge_0_avalon_master_writedata;                                           // i2c_cont_bridge_0:mstr_data_out -> i2c_cont_bridge_0_avalon_master_translator:av_writedata
	wire   [9:0] i2c_cont_bridge_0_avalon_master_address;                                             // i2c_cont_bridge_0:mstr_address -> i2c_cont_bridge_0_avalon_master_translator:av_address
	wire         i2c_cont_bridge_0_avalon_master_chipselect;                                          // i2c_cont_bridge_0:mstr_en_n -> i2c_cont_bridge_0_avalon_master_translator:av_chipselect
	wire         i2c_cont_bridge_0_avalon_master_write;                                               // i2c_cont_bridge_0:mstr_write_n -> i2c_cont_bridge_0_avalon_master_translator:av_write
	wire         i2c_cont_bridge_0_avalon_master_read;                                                // i2c_cont_bridge_0:mstr_read_n -> i2c_cont_bridge_0_avalon_master_translator:av_read
	wire  [31:0] i2c_cont_bridge_0_avalon_master_readdata;                                            // i2c_cont_bridge_0_avalon_master_translator:av_readdata -> i2c_cont_bridge_0:mstr_data_in
	wire         i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest;    // opencores_i2c_0_avalon_slave_0_translator:uav_waitrequest -> i2c_cont_bridge_0_avalon_master_translator:uav_waitrequest
	wire   [2:0] i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount;     // i2c_cont_bridge_0_avalon_master_translator:uav_burstcount -> opencores_i2c_0_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_writedata;      // i2c_cont_bridge_0_avalon_master_translator:uav_writedata -> opencores_i2c_0_avalon_slave_0_translator:uav_writedata
	wire   [9:0] i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_address;        // i2c_cont_bridge_0_avalon_master_translator:uav_address -> opencores_i2c_0_avalon_slave_0_translator:uav_address
	wire         i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_lock;           // i2c_cont_bridge_0_avalon_master_translator:uav_lock -> opencores_i2c_0_avalon_slave_0_translator:uav_lock
	wire         i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_write;          // i2c_cont_bridge_0_avalon_master_translator:uav_write -> opencores_i2c_0_avalon_slave_0_translator:uav_write
	wire         i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_read;           // i2c_cont_bridge_0_avalon_master_translator:uav_read -> opencores_i2c_0_avalon_slave_0_translator:uav_read
	wire  [31:0] i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_readdata;       // opencores_i2c_0_avalon_slave_0_translator:uav_readdata -> i2c_cont_bridge_0_avalon_master_translator:uav_readdata
	wire         i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess;    // i2c_cont_bridge_0_avalon_master_translator:uav_debugaccess -> opencores_i2c_0_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable;     // i2c_cont_bridge_0_avalon_master_translator:uav_byteenable -> opencores_i2c_0_avalon_slave_0_translator:uav_byteenable
	wire         i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid;  // opencores_i2c_0_avalon_slave_0_translator:uav_readdatavalid -> i2c_cont_bridge_0_avalon_master_translator:uav_readdatavalid
	wire         opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest;           // opencores_i2c_0:wb_ack_o -> opencores_i2c_0_avalon_slave_0_translator:av_waitrequest
	wire   [7:0] opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;             // opencores_i2c_0_avalon_slave_0_translator:av_writedata -> opencores_i2c_0:wb_dat_i
	wire   [2:0] opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_address;               // opencores_i2c_0_avalon_slave_0_translator:av_address -> opencores_i2c_0:wb_adr_i
	wire         opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;            // opencores_i2c_0_avalon_slave_0_translator:av_chipselect -> opencores_i2c_0:wb_stb_i
	wire         opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                 // opencores_i2c_0_avalon_slave_0_translator:av_write -> opencores_i2c_0:wb_we_i
	wire   [7:0] opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;              // opencores_i2c_0:wb_dat_o -> opencores_i2c_0_avalon_slave_0_translator:av_readdata
	wire         rst_controller_reset_out_reset;                                                      // rst_controller:reset_out -> [i2c_cont_bridge_0:reset_n, i2c_cont_bridge_0_avalon_master_translator:reset, i2c_cont_bridge_0_slv_translator:reset, opencores_i2c_0:wb_rst_i, opencores_i2c_0_avalon_slave_0_translator:reset, vj_avalon_master_0:reset_n, vj_avalon_master_0_avalon_master_translator:reset]

	vj_avalon_master vj_avalon_master_0 (
		.clk           (clk_clk),                                       //       clock_sink.clk
		.reset_n       (~rst_controller_reset_out_reset),               // clock_sink_reset.reset_n
		.read_n        (vj_avalon_master_0_avalon_master_read),         //    avalon_master.read_n
		.write_n       (vj_avalon_master_0_avalon_master_write),        //                 .write_n
		.address       (vj_avalon_master_0_avalon_master_address),      //                 .address
		.data_out      (vj_avalon_master_0_avalon_master_writedata),    //                 .writedata
		.waitrequest_n (~vj_avalon_master_0_avalon_master_waitrequest), //                 .waitrequest_n
		.data_in       (vj_avalon_master_0_avalon_master_readdata),     //                 .readdata
		.clk_pls_p     (vj_clk_pls_p_export)                            //        clk_pls_p.export
	);

	i2c_cont_bridge i2c_cont_bridge_0 (
		.reset_n            (~rst_controller_reset_out_reset),                                  //         reset.reset_n
		.clk                (clk_clk),                                                          //         clock.clk
		.slv_address        (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_address),     //           slv.address
		.slv_read_n         (~i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_read),       //              .read_n
		.slv_write_n        (~i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_write),      //              .write_n
		.slv_data_in        (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_writedata),   //              .writedata
		.slv_waitrequest_n  (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_waitrequest), //              .waitrequest_n
		.slv_data_out       (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_readdata),    //              .readdata
		.slv_en_n           (~i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_chipselect), //              .chipselect_n
		.mstr_en_n          (i2c_cont_bridge_0_avalon_master_chipselect),                       // avalon_master.chipselect_n
		.mstr_address       (i2c_cont_bridge_0_avalon_master_address),                          //              .address
		.mstr_write_n       (i2c_cont_bridge_0_avalon_master_write),                            //              .write_n
		.mstr_read_n        (i2c_cont_bridge_0_avalon_master_read),                             //              .read_n
		.mstr_data_in       (i2c_cont_bridge_0_avalon_master_readdata),                         //              .readdata
		.mstr_data_out      (i2c_cont_bridge_0_avalon_master_writedata),                        //              .writedata
		.mstr_waitrequest_n (~i2c_cont_bridge_0_avalon_master_waitrequest)                      //              .waitrequest_n
	);

	opencores_i2c opencores_i2c_0 (
		.wb_clk_i   (clk_clk),                                                                   //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                            //      clock_reset.reset
		.scl_pad_io (opencores_i2c_0_export_0_scl_pad_io),                                       //         export_0.export
		.sda_pad_io (opencores_i2c_0_export_0_sda_pad_io),                                       //                 .export
		.wb_adr_i   (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                 .readdata
		.wb_we_i    (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_write),       //                 .write
		.wb_stb_i   (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  ()                                                                           // interrupt_sender.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) vj_avalon_master_0_avalon_master_translator (
		.clk                   (clk_clk),                                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                     reset.reset
		.uav_address           (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (vj_avalon_master_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (vj_avalon_master_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_read               (~vj_avalon_master_0_avalon_master_read),                                              //                          .read
		.av_readdata           (vj_avalon_master_0_avalon_master_readdata),                                           //                          .readdata
		.av_write              (~vj_avalon_master_0_avalon_master_write),                                             //                          .write
		.av_writedata          (vj_avalon_master_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                                //               (terminated)
		.av_byteenable         (4'b1111),                                                                             //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                                //               (terminated)
		.av_chipselect         (1'b0),                                                                                //               (terminated)
		.av_readdatavalid      (),                                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                                //               (terminated)
		.av_debugaccess        (1'b0),                                                                                //               (terminated)
		.uav_clken             (),                                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                                 //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_cont_bridge_0_slv_translator (
		.clk                   (clk_clk),                                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (vj_avalon_master_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_address),                        //      avalon_anti_slave_0.address
		.av_write              (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_write),                          //                         .write
		.av_read               (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_read),                           //                         .read
		.av_readdata           (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_readdata),                       //                         .readdata
		.av_writedata          (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_writedata),                      //                         .writedata
		.av_waitrequest        (~i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_waitrequest),                   //                         .waitrequest
		.av_chipselect         (i2c_cont_bridge_0_slv_translator_avalon_anti_slave_0_chipselect),                     //                         .chipselect
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) i2c_cont_bridge_0_avalon_master_translator (
		.clk                   (clk_clk),                                                                            //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address           (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (i2c_cont_bridge_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (i2c_cont_bridge_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_chipselect         (~i2c_cont_bridge_0_avalon_master_chipselect),                                        //                          .chipselect
		.av_read               (~i2c_cont_bridge_0_avalon_master_read),                                              //                          .read
		.av_readdata           (i2c_cont_bridge_0_avalon_master_readdata),                                           //                          .readdata
		.av_write              (~i2c_cont_bridge_0_avalon_master_write),                                             //                          .write
		.av_writedata          (i2c_cont_bridge_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_readdatavalid      (),                                                                                   //               (terminated)
		.av_lock               (1'b0),                                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) opencores_i2c_0_avalon_slave_0_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (i2c_cont_bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address            (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_address),              //      avalon_anti_slave_0.address
		.av_write              (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                //                         .write
		.av_readdata           (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),             //                         .readdata
		.av_writedata          (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),            //                         .writedata
		.av_waitrequest        (~opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest),         //                         .waitrequest
		.av_chipselect         (opencores_i2c_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),           //                         .chipselect
		.av_read               (),                                                                                   //              (terminated)
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
